// moore state machine
// 9 states
// 1 input
// 1 output

module ();
endmodule